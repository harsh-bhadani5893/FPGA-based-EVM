library verilog;
use verilog.vl_types.all;
entity EVM_tb is
end EVM_tb;
